module top(
	input ck,reset,
	output [7:0]red,green,
	output [7:0]ctrl
);



endmodule
